MYCIRCUIT.CIR
T1      1       4       2       4       Z0=3.34893107629129 F=1.0 NL=0.125
T2      2       5       0       6       Z0=1.4051505242882971 F=1.0 NL=0.125
T3      2       7       3       7       Z0=3.3489310762912896 F=1.0 NL=0.125
.END
