MYCIRCUIT.CIR
L1          1           2           3.34893107629129
C2          2           0           0.711667527937262
L3          2           3           3.3489310762912896
.END
