MYCIRCUIT.CIR
T1      1       2       4       4       Z0=3.3489310762912896 F=1.0 NL=0.125
T2      2       0       5       6       Z0=1.405150524288297 F=1.0 NL=0.125
T3      2       3       7       7       Z0=3.348931076291289 F=1.0 NL=0.125
.END
